// pcihellocore.v

// Generated using ACDS version 12.1 177 at 2013.06.18.08:24:05

`timescale 1 ps / 1 ps
module pcihellocore (
		input  wire        pcie_hard_ip_0_powerdown_pll_powerdown, //    pcie_hard_ip_0_powerdown.pll_powerdown
		input  wire        pcie_hard_ip_0_powerdown_gxb_powerdown, //                            .gxb_powerdown
		output wire        pcie_hard_ip_0_tx_out_tx_dataout_0,     //       pcie_hard_ip_0_tx_out.tx_dataout_0
		output wire [31:0] hexport_external_connection_export,     // hexport_external_connection.export
		input  wire [15:0] inport_external_connection_export,      //  inport_external_connection.export
		input  wire        pcie_hard_ip_0_pcie_rstn_export,        //    pcie_hard_ip_0_pcie_rstn.export
		input  wire        pcie_hard_ip_0_refclk_export,           //       pcie_hard_ip_0_refclk.export
		input  wire        pcie_hard_ip_0_rx_in_rx_datain_0        //        pcie_hard_ip_0_rx_in.rx_datain_0
	);

	wire          pcie_hard_ip_0_pcie_core_clk_clk;                                                        // pcie_hard_ip_0:pcie_core_clk_clk -> [addr_router:clk, burst_adapter:clk, burst_adapter_001:clk, burst_adapter_002:clk, cmd_xbar_demux:clk, hexport:clk, hexport_s1_translator:clk, hexport_s1_translator_avalon_universal_slave_0_agent:clk, hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, id_router:clk, id_router_001:clk, id_router_002:clk, id_router_003:clk, inport:clk, inport_s1_translator:clk, inport_s1_translator_avalon_universal_slave_0_agent:clk, inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, irq_mapper:clk, irq_synchronizer:receiver_clk, irq_synchronizer:sender_clk, limiter:clk, pcie_hard_ip_0:cal_blk_clk_clk, pcie_hard_ip_0:fixedclk_clk, pcie_hard_ip_0:reconfig_gxbclk_clk, pcie_hard_ip_0_bar0_translator:clk, pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:clk, pcie_hard_ip_0_cra_translator:clk, pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:clk, pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, pcie_hard_ip_0_txs_translator:clk, pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:clk, pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, rsp_xbar_demux:clk, rsp_xbar_demux_001:clk, rsp_xbar_demux_002:clk, rsp_xbar_demux_003:clk, rsp_xbar_mux:clk, rst_controller:clk, width_adapter:clk, width_adapter_001:clk, width_adapter_002:clk, width_adapter_003:clk, width_adapter_004:clk, width_adapter_005:clk]
	wire    [6:0] pcie_hard_ip_0_bar0_burstcount;                                                          // pcie_hard_ip_0:bar0_burstcount -> pcie_hard_ip_0_bar0_translator:av_burstcount
	wire          pcie_hard_ip_0_bar0_waitrequest;                                                         // pcie_hard_ip_0_bar0_translator:av_waitrequest -> pcie_hard_ip_0:bar0_waitrequest
	wire   [63:0] pcie_hard_ip_0_bar0_writedata;                                                           // pcie_hard_ip_0:bar0_writedata -> pcie_hard_ip_0_bar0_translator:av_writedata
	wire   [31:0] pcie_hard_ip_0_bar0_address;                                                             // pcie_hard_ip_0:bar0_address -> pcie_hard_ip_0_bar0_translator:av_address
	wire          pcie_hard_ip_0_bar0_write;                                                               // pcie_hard_ip_0:bar0_write -> pcie_hard_ip_0_bar0_translator:av_write
	wire          pcie_hard_ip_0_bar0_read;                                                                // pcie_hard_ip_0:bar0_read -> pcie_hard_ip_0_bar0_translator:av_read
	wire   [63:0] pcie_hard_ip_0_bar0_readdata;                                                            // pcie_hard_ip_0_bar0_translator:av_readdata -> pcie_hard_ip_0:bar0_readdata
	wire    [7:0] pcie_hard_ip_0_bar0_byteenable;                                                          // pcie_hard_ip_0:bar0_byteenable -> pcie_hard_ip_0_bar0_translator:av_byteenable
	wire          pcie_hard_ip_0_bar0_readdatavalid;                                                       // pcie_hard_ip_0_bar0_translator:av_readdatavalid -> pcie_hard_ip_0:bar0_readdatavalid
	wire          pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_waitrequest;                           // pcie_hard_ip_0:cra_waitrequest -> pcie_hard_ip_0_cra_translator:av_waitrequest
	wire   [31:0] pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_writedata;                             // pcie_hard_ip_0_cra_translator:av_writedata -> pcie_hard_ip_0:cra_writedata
	wire   [11:0] pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_address;                               // pcie_hard_ip_0_cra_translator:av_address -> pcie_hard_ip_0:cra_address
	wire          pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_chipselect;                            // pcie_hard_ip_0_cra_translator:av_chipselect -> pcie_hard_ip_0:cra_chipselect
	wire          pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_write;                                 // pcie_hard_ip_0_cra_translator:av_write -> pcie_hard_ip_0:cra_write
	wire          pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_read;                                  // pcie_hard_ip_0_cra_translator:av_read -> pcie_hard_ip_0:cra_read
	wire   [31:0] pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_readdata;                              // pcie_hard_ip_0:cra_readdata -> pcie_hard_ip_0_cra_translator:av_readdata
	wire    [3:0] pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_byteenable;                            // pcie_hard_ip_0_cra_translator:av_byteenable -> pcie_hard_ip_0:cra_byteenable
	wire    [1:0] inport_s1_translator_avalon_anti_slave_0_address;                                        // inport_s1_translator:av_address -> inport:address
	wire   [31:0] inport_s1_translator_avalon_anti_slave_0_readdata;                                       // inport:readdata -> inport_s1_translator:av_readdata
	wire   [31:0] hexport_s1_translator_avalon_anti_slave_0_writedata;                                     // hexport_s1_translator:av_writedata -> hexport:writedata
	wire    [1:0] hexport_s1_translator_avalon_anti_slave_0_address;                                       // hexport_s1_translator:av_address -> hexport:address
	wire          hexport_s1_translator_avalon_anti_slave_0_chipselect;                                    // hexport_s1_translator:av_chipselect -> hexport:chipselect
	wire          hexport_s1_translator_avalon_anti_slave_0_write;                                         // hexport_s1_translator:av_write -> hexport:write_n
	wire   [31:0] hexport_s1_translator_avalon_anti_slave_0_readdata;                                      // hexport:readdata -> hexport_s1_translator:av_readdata
	wire          pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_waitrequest;                           // pcie_hard_ip_0:txs_waitrequest -> pcie_hard_ip_0_txs_translator:av_waitrequest
	wire    [6:0] pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_burstcount;                            // pcie_hard_ip_0_txs_translator:av_burstcount -> pcie_hard_ip_0:txs_burstcount
	wire   [63:0] pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_writedata;                             // pcie_hard_ip_0_txs_translator:av_writedata -> pcie_hard_ip_0:txs_writedata
	wire   [14:0] pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_address;                               // pcie_hard_ip_0_txs_translator:av_address -> pcie_hard_ip_0:txs_address
	wire          pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_chipselect;                            // pcie_hard_ip_0_txs_translator:av_chipselect -> pcie_hard_ip_0:txs_chipselect
	wire          pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_write;                                 // pcie_hard_ip_0_txs_translator:av_write -> pcie_hard_ip_0:txs_write
	wire          pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_read;                                  // pcie_hard_ip_0_txs_translator:av_read -> pcie_hard_ip_0:txs_read
	wire   [63:0] pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_readdata;                              // pcie_hard_ip_0:txs_readdata -> pcie_hard_ip_0_txs_translator:av_readdata
	wire          pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_readdatavalid;                         // pcie_hard_ip_0:txs_readdatavalid -> pcie_hard_ip_0_txs_translator:av_readdatavalid
	wire    [7:0] pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_byteenable;                            // pcie_hard_ip_0_txs_translator:av_byteenable -> pcie_hard_ip_0:txs_byteenable
	wire          pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_waitrequest;                    // pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:av_waitrequest -> pcie_hard_ip_0_bar0_translator:uav_waitrequest
	wire    [9:0] pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_burstcount;                     // pcie_hard_ip_0_bar0_translator:uav_burstcount -> pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [63:0] pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_writedata;                      // pcie_hard_ip_0_bar0_translator:uav_writedata -> pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_address;                        // pcie_hard_ip_0_bar0_translator:uav_address -> pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:av_address
	wire          pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_lock;                           // pcie_hard_ip_0_bar0_translator:uav_lock -> pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:av_lock
	wire          pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_write;                          // pcie_hard_ip_0_bar0_translator:uav_write -> pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:av_write
	wire          pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_read;                           // pcie_hard_ip_0_bar0_translator:uav_read -> pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:av_read
	wire   [63:0] pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_readdata;                       // pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:av_readdata -> pcie_hard_ip_0_bar0_translator:uav_readdata
	wire          pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_debugaccess;                    // pcie_hard_ip_0_bar0_translator:uav_debugaccess -> pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [7:0] pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_byteenable;                     // pcie_hard_ip_0_bar0_translator:uav_byteenable -> pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:av_byteenable
	wire          pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_readdatavalid;                  // pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:av_readdatavalid -> pcie_hard_ip_0_bar0_translator:uav_readdatavalid
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // pcie_hard_ip_0_cra_translator:uav_waitrequest -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_burstcount;              // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:m0_burstcount -> pcie_hard_ip_0_cra_translator:uav_burstcount
	wire   [31:0] pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_writedata;               // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:m0_writedata -> pcie_hard_ip_0_cra_translator:uav_writedata
	wire   [31:0] pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_address;                 // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:m0_address -> pcie_hard_ip_0_cra_translator:uav_address
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_write;                   // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:m0_write -> pcie_hard_ip_0_cra_translator:uav_write
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_lock;                    // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:m0_lock -> pcie_hard_ip_0_cra_translator:uav_lock
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_read;                    // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:m0_read -> pcie_hard_ip_0_cra_translator:uav_read
	wire   [31:0] pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_readdata;                // pcie_hard_ip_0_cra_translator:uav_readdata -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // pcie_hard_ip_0_cra_translator:uav_readdatavalid -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pcie_hard_ip_0_cra_translator:uav_debugaccess
	wire    [3:0] pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_byteenable;              // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:m0_byteenable -> pcie_hard_ip_0_cra_translator:uav_byteenable
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rf_source_valid;            // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rf_source_valid -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [117:0] pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rf_source_data;             // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rf_source_data -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rf_source_ready;            // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [117:0] pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          inport_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // inport_s1_translator:uav_waitrequest -> inport_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] inport_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // inport_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> inport_s1_translator:uav_burstcount
	wire   [31:0] inport_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                        // inport_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> inport_s1_translator:uav_writedata
	wire   [31:0] inport_s1_translator_avalon_universal_slave_0_agent_m0_address;                          // inport_s1_translator_avalon_universal_slave_0_agent:m0_address -> inport_s1_translator:uav_address
	wire          inport_s1_translator_avalon_universal_slave_0_agent_m0_write;                            // inport_s1_translator_avalon_universal_slave_0_agent:m0_write -> inport_s1_translator:uav_write
	wire          inport_s1_translator_avalon_universal_slave_0_agent_m0_lock;                             // inport_s1_translator_avalon_universal_slave_0_agent:m0_lock -> inport_s1_translator:uav_lock
	wire          inport_s1_translator_avalon_universal_slave_0_agent_m0_read;                             // inport_s1_translator_avalon_universal_slave_0_agent:m0_read -> inport_s1_translator:uav_read
	wire   [31:0] inport_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                         // inport_s1_translator:uav_readdata -> inport_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          inport_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // inport_s1_translator:uav_readdatavalid -> inport_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          inport_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // inport_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> inport_s1_translator:uav_debugaccess
	wire    [3:0] inport_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // inport_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> inport_s1_translator:uav_byteenable
	wire          inport_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // inport_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          inport_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // inport_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          inport_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // inport_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [117:0] inport_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                      // inport_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          inport_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> inport_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> inport_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> inport_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> inport_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [117:0] inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> inport_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // inport_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          inport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // inport_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> inport_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] inport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // inport_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> inport_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          inport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // inport_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> inport_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                     // hexport_s1_translator:uav_waitrequest -> hexport_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] hexport_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                      // hexport_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> hexport_s1_translator:uav_burstcount
	wire   [31:0] hexport_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                       // hexport_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> hexport_s1_translator:uav_writedata
	wire   [31:0] hexport_s1_translator_avalon_universal_slave_0_agent_m0_address;                         // hexport_s1_translator_avalon_universal_slave_0_agent:m0_address -> hexport_s1_translator:uav_address
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_m0_write;                           // hexport_s1_translator_avalon_universal_slave_0_agent:m0_write -> hexport_s1_translator:uav_write
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_m0_lock;                            // hexport_s1_translator_avalon_universal_slave_0_agent:m0_lock -> hexport_s1_translator:uav_lock
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_m0_read;                            // hexport_s1_translator_avalon_universal_slave_0_agent:m0_read -> hexport_s1_translator:uav_read
	wire   [31:0] hexport_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                        // hexport_s1_translator:uav_readdata -> hexport_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                   // hexport_s1_translator:uav_readdatavalid -> hexport_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                     // hexport_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> hexport_s1_translator:uav_debugaccess
	wire    [3:0] hexport_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                      // hexport_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> hexport_s1_translator:uav_byteenable
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;              // hexport_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                    // hexport_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;            // hexport_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [117:0] hexport_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                     // hexport_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                    // hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> hexport_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;           // hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> hexport_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                 // hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> hexport_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;         // hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> hexport_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [117:0] hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                  // hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> hexport_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                 // hexport_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;               // hexport_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> hexport_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [31:0] hexport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                // hexport_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> hexport_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;               // hexport_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> hexport_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // pcie_hard_ip_0_txs_translator:uav_waitrequest -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [9:0] pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_burstcount;              // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:m0_burstcount -> pcie_hard_ip_0_txs_translator:uav_burstcount
	wire   [63:0] pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_writedata;               // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:m0_writedata -> pcie_hard_ip_0_txs_translator:uav_writedata
	wire   [31:0] pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_address;                 // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:m0_address -> pcie_hard_ip_0_txs_translator:uav_address
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_write;                   // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:m0_write -> pcie_hard_ip_0_txs_translator:uav_write
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_lock;                    // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:m0_lock -> pcie_hard_ip_0_txs_translator:uav_lock
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_read;                    // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:m0_read -> pcie_hard_ip_0_txs_translator:uav_read
	wire   [63:0] pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_readdata;                // pcie_hard_ip_0_txs_translator:uav_readdata -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // pcie_hard_ip_0_txs_translator:uav_readdatavalid -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:m0_debugaccess -> pcie_hard_ip_0_txs_translator:uav_debugaccess
	wire    [7:0] pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_byteenable;              // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:m0_byteenable -> pcie_hard_ip_0_txs_translator:uav_byteenable
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rf_source_valid;            // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rf_source_valid -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [153:0] pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rf_source_data;             // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rf_source_data -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rf_source_ready;            // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [153:0] pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rf_sink_ready -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [63:0] pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent_cp_endofpacket;           // pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent_cp_valid;                 // pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent_cp_startofpacket;         // pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [152:0] pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent_cp_data;                  // pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent_cp_ready;                 // addr_router:sink_ready -> pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:cp_ready
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router:sink_endofpacket
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rp_valid;                   // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rp_valid -> id_router:sink_valid
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router:sink_startofpacket
	wire  [116:0] pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rp_data;                    // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rp_data -> id_router:sink_data
	wire          pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router:sink_ready -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:rp_ready
	wire          inport_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // inport_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_001:sink_endofpacket
	wire          inport_s1_translator_avalon_universal_slave_0_agent_rp_valid;                            // inport_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_001:sink_valid
	wire          inport_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // inport_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [116:0] inport_s1_translator_avalon_universal_slave_0_agent_rp_data;                             // inport_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_001:sink_data
	wire          inport_s1_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_001:sink_ready -> inport_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                     // hexport_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_rp_valid;                           // hexport_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                   // hexport_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [116:0] hexport_s1_translator_avalon_universal_slave_0_agent_rp_data;                            // hexport_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          hexport_s1_translator_avalon_universal_slave_0_agent_rp_ready;                           // id_router_002:sink_ready -> hexport_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rp_valid;                   // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [152:0] pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rp_data;                    // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_003:sink_ready -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                             // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                   // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                           // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [152:0] addr_router_src_data;                                                                    // addr_router:src_data -> limiter:cmd_sink_data
	wire    [3:0] addr_router_src_channel;                                                                 // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                   // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                             // limiter:rsp_src_endofpacket -> pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                   // limiter:rsp_src_valid -> pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                           // limiter:rsp_src_startofpacket -> pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [152:0] limiter_rsp_src_data;                                                                    // limiter:rsp_src_data -> pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:rp_data
	wire    [3:0] limiter_rsp_src_channel;                                                                 // limiter:rsp_src_channel -> pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                   // pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                       // burst_adapter:source0_endofpacket -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                             // burst_adapter:source0_valid -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                     // burst_adapter:source0_startofpacket -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [116:0] burst_adapter_source0_data;                                                              // burst_adapter:source0_data -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                             // pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire    [3:0] burst_adapter_source0_channel;                                                           // burst_adapter:source0_channel -> pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                   // burst_adapter_001:source0_endofpacket -> inport_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                         // burst_adapter_001:source0_valid -> inport_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                 // burst_adapter_001:source0_startofpacket -> inport_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [116:0] burst_adapter_001_source0_data;                                                          // burst_adapter_001:source0_data -> inport_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                         // inport_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire    [3:0] burst_adapter_001_source0_channel;                                                       // burst_adapter_001:source0_channel -> inport_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_002_source0_endofpacket;                                                   // burst_adapter_002:source0_endofpacket -> hexport_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_002_source0_valid;                                                         // burst_adapter_002:source0_valid -> hexport_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_002_source0_startofpacket;                                                 // burst_adapter_002:source0_startofpacket -> hexport_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [116:0] burst_adapter_002_source0_data;                                                          // burst_adapter_002:source0_data -> hexport_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_002_source0_ready;                                                         // hexport_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire    [3:0] burst_adapter_002_source0_channel;                                                       // burst_adapter_002:source0_channel -> hexport_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rst_controller_reset_out_reset;                                                          // rst_controller:reset_out -> [addr_router:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, cmd_xbar_demux:reset, hexport:reset_n, hexport_s1_translator:reset, hexport_s1_translator_avalon_universal_slave_0_agent:reset, hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router:reset, id_router_001:reset, id_router_002:reset, id_router_003:reset, inport:reset_n, inport_s1_translator:reset, inport_s1_translator_avalon_universal_slave_0_agent:reset, inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, pcie_hard_ip_0_bar0_translator:reset, pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent:reset, pcie_hard_ip_0_cra_translator:reset, pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent:reset, pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pcie_hard_ip_0_txs_translator:reset, pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:reset, pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_mux:reset, width_adapter:reset, width_adapter_001:reset, width_adapter_002:reset, width_adapter_003:reset, width_adapter_004:reset, width_adapter_005:reset]
	wire          pcie_hard_ip_0_pcie_core_reset_reset;                                                    // pcie_hard_ip_0:pcie_core_reset_reset_n -> [irq_mapper:reset, irq_synchronizer:receiver_reset, irq_synchronizer:sender_reset, rst_controller:reset_in0]
	wire          cmd_xbar_demux_src0_endofpacket;                                                         // cmd_xbar_demux:src0_endofpacket -> width_adapter:in_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                               // cmd_xbar_demux:src0_valid -> width_adapter:in_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                       // cmd_xbar_demux:src0_startofpacket -> width_adapter:in_startofpacket
	wire  [152:0] cmd_xbar_demux_src0_data;                                                                // cmd_xbar_demux:src0_data -> width_adapter:in_data
	wire    [3:0] cmd_xbar_demux_src0_channel;                                                             // cmd_xbar_demux:src0_channel -> width_adapter:in_channel
	wire          cmd_xbar_demux_src1_endofpacket;                                                         // cmd_xbar_demux:src1_endofpacket -> width_adapter_002:in_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                               // cmd_xbar_demux:src1_valid -> width_adapter_002:in_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                       // cmd_xbar_demux:src1_startofpacket -> width_adapter_002:in_startofpacket
	wire  [152:0] cmd_xbar_demux_src1_data;                                                                // cmd_xbar_demux:src1_data -> width_adapter_002:in_data
	wire    [3:0] cmd_xbar_demux_src1_channel;                                                             // cmd_xbar_demux:src1_channel -> width_adapter_002:in_channel
	wire          cmd_xbar_demux_src2_endofpacket;                                                         // cmd_xbar_demux:src2_endofpacket -> width_adapter_004:in_endofpacket
	wire          cmd_xbar_demux_src2_valid;                                                               // cmd_xbar_demux:src2_valid -> width_adapter_004:in_valid
	wire          cmd_xbar_demux_src2_startofpacket;                                                       // cmd_xbar_demux:src2_startofpacket -> width_adapter_004:in_startofpacket
	wire  [152:0] cmd_xbar_demux_src2_data;                                                                // cmd_xbar_demux:src2_data -> width_adapter_004:in_data
	wire    [3:0] cmd_xbar_demux_src2_channel;                                                             // cmd_xbar_demux:src2_channel -> width_adapter_004:in_channel
	wire          cmd_xbar_demux_src3_endofpacket;                                                         // cmd_xbar_demux:src3_endofpacket -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          cmd_xbar_demux_src3_valid;                                                               // cmd_xbar_demux:src3_valid -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:cp_valid
	wire          cmd_xbar_demux_src3_startofpacket;                                                       // cmd_xbar_demux:src3_startofpacket -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [152:0] cmd_xbar_demux_src3_data;                                                                // cmd_xbar_demux:src3_data -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:cp_data
	wire    [3:0] cmd_xbar_demux_src3_channel;                                                             // cmd_xbar_demux:src3_channel -> pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:cp_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                         // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                               // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                       // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [152:0] rsp_xbar_demux_src0_data;                                                                // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire    [3:0] rsp_xbar_demux_src0_channel;                                                             // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                               // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                     // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                           // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                   // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [152:0] rsp_xbar_demux_001_src0_data;                                                            // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire    [3:0] rsp_xbar_demux_001_src0_channel;                                                         // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                           // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                     // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux:sink2_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                           // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux:sink2_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                   // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux:sink2_startofpacket
	wire  [152:0] rsp_xbar_demux_002_src0_data;                                                            // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux:sink2_data
	wire    [3:0] rsp_xbar_demux_002_src0_channel;                                                         // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux:sink2_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                           // rsp_xbar_mux:sink2_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                     // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux:sink3_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                           // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux:sink3_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                   // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux:sink3_startofpacket
	wire  [152:0] rsp_xbar_demux_003_src0_data;                                                            // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux:sink3_data
	wire    [3:0] rsp_xbar_demux_003_src0_channel;                                                         // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux:sink3_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                           // rsp_xbar_mux:sink3_ready -> rsp_xbar_demux_003:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                             // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                           // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [152:0] limiter_cmd_src_data;                                                                    // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire    [3:0] limiter_cmd_src_channel;                                                                 // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                   // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                            // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                  // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                          // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [152:0] rsp_xbar_mux_src_data;                                                                   // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire    [3:0] rsp_xbar_mux_src_channel;                                                                // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                  // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          cmd_xbar_demux_src3_ready;                                                               // pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent:cp_ready -> cmd_xbar_demux:src3_ready
	wire          id_router_003_src_endofpacket;                                                           // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                 // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                         // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [152:0] id_router_003_src_data;                                                                  // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [3:0] id_router_003_src_channel;                                                               // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                 // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_demux_src0_ready;                                                               // width_adapter:in_ready -> cmd_xbar_demux:src0_ready
	wire          width_adapter_src_endofpacket;                                                           // width_adapter:out_endofpacket -> burst_adapter:sink0_endofpacket
	wire          width_adapter_src_valid;                                                                 // width_adapter:out_valid -> burst_adapter:sink0_valid
	wire          width_adapter_src_startofpacket;                                                         // width_adapter:out_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [116:0] width_adapter_src_data;                                                                  // width_adapter:out_data -> burst_adapter:sink0_data
	wire          width_adapter_src_ready;                                                                 // burst_adapter:sink0_ready -> width_adapter:out_ready
	wire    [3:0] width_adapter_src_channel;                                                               // width_adapter:out_channel -> burst_adapter:sink0_channel
	wire          id_router_src_endofpacket;                                                               // id_router:src_endofpacket -> width_adapter_001:in_endofpacket
	wire          id_router_src_valid;                                                                     // id_router:src_valid -> width_adapter_001:in_valid
	wire          id_router_src_startofpacket;                                                             // id_router:src_startofpacket -> width_adapter_001:in_startofpacket
	wire  [116:0] id_router_src_data;                                                                      // id_router:src_data -> width_adapter_001:in_data
	wire    [3:0] id_router_src_channel;                                                                   // id_router:src_channel -> width_adapter_001:in_channel
	wire          id_router_src_ready;                                                                     // width_adapter_001:in_ready -> id_router:src_ready
	wire          width_adapter_001_src_endofpacket;                                                       // width_adapter_001:out_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          width_adapter_001_src_valid;                                                             // width_adapter_001:out_valid -> rsp_xbar_demux:sink_valid
	wire          width_adapter_001_src_startofpacket;                                                     // width_adapter_001:out_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [152:0] width_adapter_001_src_data;                                                              // width_adapter_001:out_data -> rsp_xbar_demux:sink_data
	wire          width_adapter_001_src_ready;                                                             // rsp_xbar_demux:sink_ready -> width_adapter_001:out_ready
	wire    [3:0] width_adapter_001_src_channel;                                                           // width_adapter_001:out_channel -> rsp_xbar_demux:sink_channel
	wire          cmd_xbar_demux_src1_ready;                                                               // width_adapter_002:in_ready -> cmd_xbar_demux:src1_ready
	wire          width_adapter_002_src_endofpacket;                                                       // width_adapter_002:out_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          width_adapter_002_src_valid;                                                             // width_adapter_002:out_valid -> burst_adapter_001:sink0_valid
	wire          width_adapter_002_src_startofpacket;                                                     // width_adapter_002:out_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire  [116:0] width_adapter_002_src_data;                                                              // width_adapter_002:out_data -> burst_adapter_001:sink0_data
	wire          width_adapter_002_src_ready;                                                             // burst_adapter_001:sink0_ready -> width_adapter_002:out_ready
	wire    [3:0] width_adapter_002_src_channel;                                                           // width_adapter_002:out_channel -> burst_adapter_001:sink0_channel
	wire          id_router_001_src_endofpacket;                                                           // id_router_001:src_endofpacket -> width_adapter_003:in_endofpacket
	wire          id_router_001_src_valid;                                                                 // id_router_001:src_valid -> width_adapter_003:in_valid
	wire          id_router_001_src_startofpacket;                                                         // id_router_001:src_startofpacket -> width_adapter_003:in_startofpacket
	wire  [116:0] id_router_001_src_data;                                                                  // id_router_001:src_data -> width_adapter_003:in_data
	wire    [3:0] id_router_001_src_channel;                                                               // id_router_001:src_channel -> width_adapter_003:in_channel
	wire          id_router_001_src_ready;                                                                 // width_adapter_003:in_ready -> id_router_001:src_ready
	wire          width_adapter_003_src_endofpacket;                                                       // width_adapter_003:out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          width_adapter_003_src_valid;                                                             // width_adapter_003:out_valid -> rsp_xbar_demux_001:sink_valid
	wire          width_adapter_003_src_startofpacket;                                                     // width_adapter_003:out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [152:0] width_adapter_003_src_data;                                                              // width_adapter_003:out_data -> rsp_xbar_demux_001:sink_data
	wire          width_adapter_003_src_ready;                                                             // rsp_xbar_demux_001:sink_ready -> width_adapter_003:out_ready
	wire    [3:0] width_adapter_003_src_channel;                                                           // width_adapter_003:out_channel -> rsp_xbar_demux_001:sink_channel
	wire          cmd_xbar_demux_src2_ready;                                                               // width_adapter_004:in_ready -> cmd_xbar_demux:src2_ready
	wire          width_adapter_004_src_endofpacket;                                                       // width_adapter_004:out_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire          width_adapter_004_src_valid;                                                             // width_adapter_004:out_valid -> burst_adapter_002:sink0_valid
	wire          width_adapter_004_src_startofpacket;                                                     // width_adapter_004:out_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire  [116:0] width_adapter_004_src_data;                                                              // width_adapter_004:out_data -> burst_adapter_002:sink0_data
	wire          width_adapter_004_src_ready;                                                             // burst_adapter_002:sink0_ready -> width_adapter_004:out_ready
	wire    [3:0] width_adapter_004_src_channel;                                                           // width_adapter_004:out_channel -> burst_adapter_002:sink0_channel
	wire          id_router_002_src_endofpacket;                                                           // id_router_002:src_endofpacket -> width_adapter_005:in_endofpacket
	wire          id_router_002_src_valid;                                                                 // id_router_002:src_valid -> width_adapter_005:in_valid
	wire          id_router_002_src_startofpacket;                                                         // id_router_002:src_startofpacket -> width_adapter_005:in_startofpacket
	wire  [116:0] id_router_002_src_data;                                                                  // id_router_002:src_data -> width_adapter_005:in_data
	wire    [3:0] id_router_002_src_channel;                                                               // id_router_002:src_channel -> width_adapter_005:in_channel
	wire          id_router_002_src_ready;                                                                 // width_adapter_005:in_ready -> id_router_002:src_ready
	wire          width_adapter_005_src_endofpacket;                                                       // width_adapter_005:out_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          width_adapter_005_src_valid;                                                             // width_adapter_005:out_valid -> rsp_xbar_demux_002:sink_valid
	wire          width_adapter_005_src_startofpacket;                                                     // width_adapter_005:out_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [152:0] width_adapter_005_src_data;                                                              // width_adapter_005:out_data -> rsp_xbar_demux_002:sink_data
	wire          width_adapter_005_src_ready;                                                             // rsp_xbar_demux_002:sink_ready -> width_adapter_005:out_ready
	wire    [3:0] width_adapter_005_src_channel;                                                           // width_adapter_005:out_channel -> rsp_xbar_demux_002:sink_channel
	wire    [3:0] limiter_cmd_valid_data;                                                                  // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire   [15:0] pcie_hard_ip_0_rxm_irq_irq;                                                              // irq_synchronizer:sender_irq -> pcie_hard_ip_0:rxm_irq_irq
	wire   [15:0] irq_synchronizer_receiver_irq;                                                           // irq_mapper:sender_irq -> irq_synchronizer:receiver_irq

	pcihellocore_hexport hexport (
		.clk        (pcie_hard_ip_0_pcie_core_clk_clk),                     //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (hexport_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~hexport_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (hexport_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (hexport_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (hexport_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (hexport_external_connection_export)                    // external_connection.export
	);

	pcihellocore_inport inport (
		.clk      (pcie_hard_ip_0_pcie_core_clk_clk),                  //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                   //               reset.reset_n
		.address  (inport_s1_translator_avalon_anti_slave_0_address),  //                  s1.address
		.readdata (inport_s1_translator_avalon_anti_slave_0_readdata), //                    .readdata
		.in_port  (inport_external_connection_export)                  // external_connection.export
	);

	pcihellocore_pcie_hard_ip_0 #(
		.p_pcie_hip_type                     ("2"),
		.lane_mask                           (8'b11111110),
		.max_link_width                      (1),
		.millisecond_cycle_count             ("125000"),
		.enable_gen2_core                    ("false"),
		.gen2_lane_rate_mode                 ("false"),
		.no_soft_reset                       ("false"),
		.core_clk_divider                    (2),
		.enable_ch0_pclk_out                 ("true"),
		.core_clk_source                     ("pclk"),
		.CB_P2A_AVALON_ADDR_B0               (0),
		.bar0_size_mask                      (16),
		.bar0_io_space                       ("false"),
		.bar0_64bit_mem_space                ("false"),
		.bar0_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B1               (0),
		.bar1_size_mask                      (0),
		.bar1_io_space                       ("false"),
		.bar1_64bit_mem_space                ("false"),
		.bar1_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B2               (0),
		.bar2_size_mask                      (0),
		.bar2_io_space                       ("false"),
		.bar2_64bit_mem_space                ("false"),
		.bar2_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B3               (0),
		.bar3_size_mask                      (0),
		.bar3_io_space                       ("false"),
		.bar3_64bit_mem_space                ("false"),
		.bar3_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B4               (0),
		.bar4_size_mask                      (0),
		.bar4_io_space                       ("false"),
		.bar4_64bit_mem_space                ("false"),
		.bar4_prefetchable                   ("false"),
		.CB_P2A_AVALON_ADDR_B5               (0),
		.bar5_size_mask                      (0),
		.bar5_io_space                       ("false"),
		.bar5_64bit_mem_space                ("false"),
		.bar5_prefetchable                   ("false"),
		.vendor_id                           (4466),
		.device_id                           (4),
		.revision_id                         (1),
		.class_code                          (0),
		.subsystem_vendor_id                 (4466),
		.subsystem_device_id                 (4),
		.port_link_number                    (1),
		.msi_function_count                  (0),
		.enable_msi_64bit_addressing         ("true"),
		.enable_function_msix_support        ("false"),
		.eie_before_nfts_count               (4),
		.enable_completion_timeout_disable   ("false"),
		.completion_timeout                  ("NONE"),
		.enable_adapter_half_rate_mode       ("false"),
		.msix_pba_bir                        (0),
		.msix_pba_offset                     (0),
		.msix_table_bir                      (0),
		.msix_table_offset                   (0),
		.msix_table_size                     (0),
		.use_crc_forwarding                  ("false"),
		.surprise_down_error_support         ("false"),
		.dll_active_report_support           ("false"),
		.bar_io_window_size                  ("32BIT"),
		.bar_prefetchable                    (32),
		.hot_plug_support                    (7'b0000000),
		.no_command_completed                ("true"),
		.slot_power_limit                    (0),
		.slot_power_scale                    (0),
		.slot_number                         (0),
		.enable_slot_register                ("false"),
		.advanced_errors                     ("false"),
		.enable_ecrc_check                   ("false"),
		.enable_ecrc_gen                     ("false"),
		.max_payload_size                    (0),
		.retry_buffer_last_active_address    (255),
		.credit_buffer_allocation_aux        ("ABSOLUTE"),
		.vc0_rx_flow_ctrl_posted_header      (28),
		.vc0_rx_flow_ctrl_posted_data        (198),
		.vc0_rx_flow_ctrl_nonposted_header   (30),
		.vc0_rx_flow_ctrl_nonposted_data     (0),
		.vc0_rx_flow_ctrl_compl_header       (48),
		.vc0_rx_flow_ctrl_compl_data         (256),
		.RX_BUF                              (9),
		.RH_NUM                              (7),
		.G_TAG_NUM0                          (32),
		.endpoint_l0_latency                 (0),
		.endpoint_l1_latency                 (0),
		.enable_l1_aspm                      ("false"),
		.l01_entry_latency                   (31),
		.diffclock_nfts_count                (255),
		.sameclock_nfts_count                (255),
		.l1_exit_latency_sameclock           (7),
		.l1_exit_latency_diffclock           (7),
		.l0_exit_latency_sameclock           (7),
		.l0_exit_latency_diffclock           (7),
		.gen2_diffclock_nfts_count           (255),
		.gen2_sameclock_nfts_count           (255),
		.CG_COMMON_CLOCK_MODE                (1),
		.CB_PCIE_MODE                        (0),
		.AST_LITE                            (0),
		.CB_PCIE_RX_LITE                     (0),
		.CG_RXM_IRQ_NUM                      (16),
		.CG_AVALON_S_ADDR_WIDTH              (20),
		.bypass_tl                           ("false"),
		.CG_IMPL_CRA_AV_SLAVE_PORT           (1),
		.CG_NO_CPL_REORDERING                (0),
		.CG_ENABLE_A2P_INTERRUPT             (0),
		.CG_IRQ_BIT_ENA                      (65535),
		.CB_A2P_ADDR_MAP_IS_FIXED            (1),
		.CB_A2P_ADDR_MAP_NUM_ENTRIES         (1),
		.CB_A2P_ADDR_MAP_PASS_THRU_BITS      (15),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_0_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_0_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_1_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_1_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_2_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_2_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_3_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_3_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_4_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_4_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_5_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_5_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_6_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_6_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_7_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_7_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_8_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_8_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_9_HIGH  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_9_LOW   (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_10_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_10_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_11_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_11_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_12_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_12_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_13_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_13_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_14_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_14_LOW  (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_15_HIGH (32'b00000000000000000000000000000000),
		.CB_A2P_ADDR_MAP_FIXED_TABLE_15_LOW  (32'b00000000000000000000000000000000),
		.RXM_DATA_WIDTH                      (64),
		.RXM_BEN_WIDTH                       (8),
		.TL_SELECTION                        (1),
		.pcie_mode                           ("SHARED_MODE"),
		.single_rx_detect                    (1),
		.enable_coreclk_out_half_rate        ("false"),
		.low_priority_vc                     (0),
		.link_width                          (1),
		.cyclone4                            (1)
	) pcie_hard_ip_0 (
		.pcie_core_clk_clk                  (pcie_hard_ip_0_pcie_core_clk_clk),                                //      pcie_core_clk.clk
		.pcie_core_reset_reset_n            (pcie_hard_ip_0_pcie_core_reset_reset),                            //    pcie_core_reset.reset_n
		.cal_blk_clk_clk                    (pcie_hard_ip_0_pcie_core_clk_clk),                                //        cal_blk_clk.clk
		.txs_address                        (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_address),       //                txs.address
		.txs_chipselect                     (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_chipselect),    //                   .chipselect
		.txs_byteenable                     (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.txs_readdata                       (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.txs_writedata                      (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.txs_read                           (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_read),          //                   .read
		.txs_write                          (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_write),         //                   .write
		.txs_burstcount                     (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_burstcount),    //                   .burstcount
		.txs_readdatavalid                  (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_readdatavalid), //                   .readdatavalid
		.txs_waitrequest                    (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_waitrequest),   //                   .waitrequest
		.refclk_export                      (pcie_hard_ip_0_refclk_export),                                    //             refclk.export
		.test_in_test_in                    (),                                                                //            test_in.test_in
		.pcie_rstn_export                   (pcie_hard_ip_0_pcie_rstn_export),                                 //          pcie_rstn.export
		.clocks_sim_clk250_export           (),                                                                //         clocks_sim.clk250_export
		.clocks_sim_clk500_export           (),                                                                //                   .clk500_export
		.clocks_sim_clk125_export           (),                                                                //                   .clk125_export
		.reconfig_busy_busy_altgxb_reconfig (),                                                                //      reconfig_busy.busy_altgxb_reconfig
		.pipe_ext_pipe_mode                 (),                                                                //           pipe_ext.pipe_mode
		.pipe_ext_phystatus_ext             (),                                                                //                   .phystatus_ext
		.pipe_ext_rate_ext                  (),                                                                //                   .rate_ext
		.pipe_ext_powerdown_ext             (),                                                                //                   .powerdown_ext
		.pipe_ext_txdetectrx_ext            (),                                                                //                   .txdetectrx_ext
		.pipe_ext_rxelecidle0_ext           (),                                                                //                   .rxelecidle0_ext
		.pipe_ext_rxdata0_ext               (),                                                                //                   .rxdata0_ext
		.pipe_ext_rxstatus0_ext             (),                                                                //                   .rxstatus0_ext
		.pipe_ext_rxvalid0_ext              (),                                                                //                   .rxvalid0_ext
		.pipe_ext_rxdatak0_ext              (),                                                                //                   .rxdatak0_ext
		.pipe_ext_txdata0_ext               (),                                                                //                   .txdata0_ext
		.pipe_ext_txdatak0_ext              (),                                                                //                   .txdatak0_ext
		.pipe_ext_rxpolarity0_ext           (),                                                                //                   .rxpolarity0_ext
		.pipe_ext_txcompl0_ext              (),                                                                //                   .txcompl0_ext
		.pipe_ext_txelecidle0_ext           (),                                                                //                   .txelecidle0_ext
		.powerdown_pll_powerdown            (pcie_hard_ip_0_powerdown_pll_powerdown),                          //          powerdown.pll_powerdown
		.powerdown_gxb_powerdown            (pcie_hard_ip_0_powerdown_gxb_powerdown),                          //                   .gxb_powerdown
		.bar0_address                       (pcie_hard_ip_0_bar0_address),                                     //               bar0.address
		.bar0_read                          (pcie_hard_ip_0_bar0_read),                                        //                   .read
		.bar0_waitrequest                   (pcie_hard_ip_0_bar0_waitrequest),                                 //                   .waitrequest
		.bar0_write                         (pcie_hard_ip_0_bar0_write),                                       //                   .write
		.bar0_readdatavalid                 (pcie_hard_ip_0_bar0_readdatavalid),                               //                   .readdatavalid
		.bar0_readdata                      (pcie_hard_ip_0_bar0_readdata),                                    //                   .readdata
		.bar0_writedata                     (pcie_hard_ip_0_bar0_writedata),                                   //                   .writedata
		.bar0_burstcount                    (pcie_hard_ip_0_bar0_burstcount),                                  //                   .burstcount
		.bar0_byteenable                    (pcie_hard_ip_0_bar0_byteenable),                                  //                   .byteenable
		.cra_chipselect                     (pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_chipselect),    //                cra.chipselect
		.cra_address                        (pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_address),       //                   .address
		.cra_byteenable                     (pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_byteenable),    //                   .byteenable
		.cra_read                           (pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_read),          //                   .read
		.cra_readdata                       (pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_readdata),      //                   .readdata
		.cra_write                          (pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_write),         //                   .write
		.cra_writedata                      (pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_writedata),     //                   .writedata
		.cra_waitrequest                    (pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_waitrequest),   //                   .waitrequest
		.cra_irq_irq                        (),                                                                //            cra_irq.irq
		.rxm_irq_irq                        (pcie_hard_ip_0_rxm_irq_irq),                                      //            rxm_irq.irq
		.rx_in_rx_datain_0                  (pcie_hard_ip_0_rx_in_rx_datain_0),                                //              rx_in.rx_datain_0
		.tx_out_tx_dataout_0                (pcie_hard_ip_0_tx_out_tx_dataout_0),                              //             tx_out.tx_dataout_0
		.reconfig_togxb_data                (),                                                                //     reconfig_togxb.data
		.reconfig_gxbclk_clk                (pcie_hard_ip_0_pcie_core_clk_clk),                                //    reconfig_gxbclk.clk
		.reconfig_fromgxb_0_data            (),                                                                // reconfig_fromgxb_0.data
		.fixedclk_clk                       (pcie_hard_ip_0_pcie_core_clk_clk)                                 //           fixedclk.clk
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (64),
		.AV_BURSTCOUNT_W             (7),
		.AV_BYTEENABLE_W             (8),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (10),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.AV_SYMBOLS_PER_WORD         (8),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) pcie_hard_ip_0_bar0_translator (
		.clk                   (pcie_hard_ip_0_pcie_core_clk_clk),                                       //                       clk.clk
		.reset                 (rst_controller_reset_out_reset),                                         //                     reset.reset
		.uav_address           (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount        (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read              (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write             (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest       (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid     (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable        (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata          (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata         (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock              (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess       (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address            (pcie_hard_ip_0_bar0_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest        (pcie_hard_ip_0_bar0_waitrequest),                                        //                          .waitrequest
		.av_burstcount         (pcie_hard_ip_0_bar0_burstcount),                                         //                          .burstcount
		.av_byteenable         (pcie_hard_ip_0_bar0_byteenable),                                         //                          .byteenable
		.av_read               (pcie_hard_ip_0_bar0_read),                                               //                          .read
		.av_readdata           (pcie_hard_ip_0_bar0_readdata),                                           //                          .readdata
		.av_readdatavalid      (pcie_hard_ip_0_bar0_readdatavalid),                                      //                          .readdatavalid
		.av_write              (pcie_hard_ip_0_bar0_write),                                              //                          .write
		.av_writedata          (pcie_hard_ip_0_bar0_writedata),                                          //                          .writedata
		.av_beginbursttransfer (1'b0),                                                                   //               (terminated)
		.av_begintransfer      (1'b0),                                                                   //               (terminated)
		.av_chipselect         (1'b0),                                                                   //               (terminated)
		.av_lock               (1'b0),                                                                   //               (terminated)
		.av_debugaccess        (1'b0),                                                                   //               (terminated)
		.uav_clken             (),                                                                       //               (terminated)
		.av_clken              (1'b1)                                                                    //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (12),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pcie_hard_ip_0_cra_translator (
		.clk                   (pcie_hard_ip_0_pcie_core_clk_clk),                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                //                    reset.reset
		.uav_address           (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable         (pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_waitrequest        (pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (pcie_hard_ip_0_cra_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_burstcount         (),                                                                              //              (terminated)
		.av_readdatavalid      (1'b0),                                                                          //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) inport_s1_translator (
		.clk                   (pcie_hard_ip_0_pcie_core_clk_clk),                                     //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                       //                    reset.reset
		.uav_address           (inport_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (inport_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (inport_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (inport_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (inport_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (inport_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (inport_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (inport_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (inport_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (inport_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (inport_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (inport_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_readdata           (inport_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_write              (),                                                                     //              (terminated)
		.av_read               (),                                                                     //              (terminated)
		.av_writedata          (),                                                                     //              (terminated)
		.av_begintransfer      (),                                                                     //              (terminated)
		.av_beginbursttransfer (),                                                                     //              (terminated)
		.av_burstcount         (),                                                                     //              (terminated)
		.av_byteenable         (),                                                                     //              (terminated)
		.av_readdatavalid      (1'b0),                                                                 //              (terminated)
		.av_waitrequest        (1'b0),                                                                 //              (terminated)
		.av_writebyteenable    (),                                                                     //              (terminated)
		.av_lock               (),                                                                     //              (terminated)
		.av_chipselect         (),                                                                     //              (terminated)
		.av_clken              (),                                                                     //              (terminated)
		.uav_clken             (1'b0),                                                                 //              (terminated)
		.av_debugaccess        (),                                                                     //              (terminated)
		.av_outputenable       ()                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) hexport_s1_translator (
		.clk                   (pcie_hard_ip_0_pcie_core_clk_clk),                                      //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address           (hexport_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (hexport_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (hexport_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (hexport_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (hexport_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (hexport_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (hexport_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (hexport_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (hexport_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (hexport_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (hexport_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (hexport_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (hexport_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata           (hexport_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (hexport_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect         (hexport_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read               (),                                                                      //              (terminated)
		.av_begintransfer      (),                                                                      //              (terminated)
		.av_beginbursttransfer (),                                                                      //              (terminated)
		.av_burstcount         (),                                                                      //              (terminated)
		.av_byteenable         (),                                                                      //              (terminated)
		.av_readdatavalid      (1'b0),                                                                  //              (terminated)
		.av_waitrequest        (1'b0),                                                                  //              (terminated)
		.av_writebyteenable    (),                                                                      //              (terminated)
		.av_lock               (),                                                                      //              (terminated)
		.av_clken              (),                                                                      //              (terminated)
		.uav_clken             (1'b0),                                                                  //              (terminated)
		.av_debugaccess        (),                                                                      //              (terminated)
		.av_outputenable       ()                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (15),
		.AV_DATA_W                      (64),
		.UAV_DATA_W                     (64),
		.AV_BURSTCOUNT_W                (7),
		.AV_BYTEENABLE_W                (8),
		.UAV_BYTEENABLE_W               (8),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (10),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.AV_SYMBOLS_PER_WORD            (8),
		.AV_ADDRESS_SYMBOLS             (1),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (1),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) pcie_hard_ip_0_txs_translator (
		.clk                   (pcie_hard_ip_0_pcie_core_clk_clk),                                              //                      clk.clk
		.reset                 (rst_controller_reset_out_reset),                                                //                    reset.reset
		.uav_address           (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount        (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read              (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write             (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest       (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid     (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable        (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata          (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata         (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock              (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess       (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address            (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write              (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read               (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata           (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata          (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_burstcount         (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_burstcount),                  //                         .burstcount
		.av_byteenable         (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid      (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest        (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect         (pcie_hard_ip_0_txs_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer      (),                                                                              //              (terminated)
		.av_beginbursttransfer (),                                                                              //              (terminated)
		.av_writebyteenable    (),                                                                              //              (terminated)
		.av_lock               (),                                                                              //              (terminated)
		.av_clken              (),                                                                              //              (terminated)
		.uav_clken             (1'b0),                                                                          //              (terminated)
		.av_debugaccess        (),                                                                              //              (terminated)
		.av_outputenable       ()                                                                               //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (146),
		.PKT_PROTECTION_L          (144),
		.PKT_BEGIN_BURST           (137),
		.PKT_BURSTWRAP_H           (129),
		.PKT_BURSTWRAP_L           (120),
		.PKT_BURST_SIZE_H          (132),
		.PKT_BURST_SIZE_L          (130),
		.PKT_BURST_TYPE_H          (134),
		.PKT_BURST_TYPE_L          (133),
		.PKT_BYTE_CNT_H            (119),
		.PKT_BYTE_CNT_L            (110),
		.PKT_ADDR_H                (103),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (104),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.PKT_TRANS_READ            (107),
		.PKT_TRANS_LOCK            (108),
		.PKT_TRANS_EXCLUSIVE       (109),
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_SRC_ID_H              (140),
		.PKT_SRC_ID_L              (139),
		.PKT_DEST_ID_H             (142),
		.PKT_DEST_ID_L             (141),
		.PKT_THREAD_ID_H           (143),
		.PKT_THREAD_ID_L           (143),
		.PKT_CACHE_H               (150),
		.PKT_CACHE_L               (147),
		.PKT_DATA_SIDEBAND_H       (136),
		.PKT_DATA_SIDEBAND_L       (136),
		.PKT_QOS_H                 (138),
		.PKT_QOS_L                 (138),
		.PKT_ADDR_SIDEBAND_H       (135),
		.PKT_ADDR_SIDEBAND_L       (135),
		.ST_DATA_W                 (153),
		.ST_CHANNEL_W              (4),
		.AV_BURSTCOUNT_W           (10),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (1023),
		.CACHE_VALUE               (4'b0000)
	) pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent (
		.clk              (pcie_hard_ip_0_pcie_core_clk_clk),                                                //       clk.clk
		.reset            (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.av_address       (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_address),                //        av.address
		.av_write         (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_write),                  //          .write
		.av_read          (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata     (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata      (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest   (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable    (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount    (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess   (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock          (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid         (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data          (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket   (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready         (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid         (limiter_rsp_src_valid),                                                           //        rp.valid
		.rp_data          (limiter_rsp_src_data),                                                            //          .data
		.rp_channel       (limiter_rsp_src_channel),                                                         //          .channel
		.rp_startofpacket (limiter_rsp_src_startofpacket),                                                   //          .startofpacket
		.rp_endofpacket   (limiter_rsp_src_endofpacket),                                                     //          .endofpacket
		.rp_ready         (limiter_rsp_src_ready)                                                            //          .ready
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (101),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (104),
		.PKT_SRC_ID_L              (103),
		.PKT_DEST_ID_H             (106),
		.PKT_DEST_ID_L             (105),
		.PKT_BURSTWRAP_H           (93),
		.PKT_BURSTWRAP_L           (84),
		.PKT_BYTE_CNT_H            (83),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (110),
		.PKT_PROTECTION_L          (108),
		.PKT_RESPONSE_STATUS_H     (116),
		.PKT_RESPONSE_STATUS_L     (115),
		.PKT_BURST_SIZE_H          (96),
		.PKT_BURST_SIZE_L          (94),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (117),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent (
		.clk                     (pcie_hard_ip_0_pcie_core_clk_clk),                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                             //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                             //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                              //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                                     //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                                       //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                           //                .channel
		.rf_sink_ready           (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (118),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pcie_hard_ip_0_pcie_core_clk_clk),                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (101),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (104),
		.PKT_SRC_ID_L              (103),
		.PKT_DEST_ID_H             (106),
		.PKT_DEST_ID_L             (105),
		.PKT_BURSTWRAP_H           (93),
		.PKT_BURSTWRAP_L           (84),
		.PKT_BYTE_CNT_H            (83),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (110),
		.PKT_PROTECTION_L          (108),
		.PKT_RESPONSE_STATUS_H     (116),
		.PKT_RESPONSE_STATUS_L     (115),
		.PKT_BURST_SIZE_H          (96),
		.PKT_BURST_SIZE_L          (94),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (117),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) inport_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pcie_hard_ip_0_pcie_core_clk_clk),                                               //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                 //       clk_reset.reset
		.m0_address              (inport_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (inport_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (inport_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (inport_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (inport_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (inport_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (inport_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (inport_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (inport_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (inport_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (inport_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (inport_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (inport_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (inport_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (inport_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (inport_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                 //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                        //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                          //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                              //                .channel
		.rf_sink_ready           (inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (inport_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (inport_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (inport_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (inport_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (inport_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (inport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (inport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (inport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (inport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (inport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (inport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (118),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pcie_hard_ip_0_pcie_core_clk_clk),                                               //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                 // clk_reset.reset
		.in_data           (inport_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (inport_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (inport_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (inport_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (inport_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (inport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                          // (terminated)
		.csr_read          (1'b0),                                                                           // (terminated)
		.csr_write         (1'b0),                                                                           // (terminated)
		.csr_readdata      (),                                                                               // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                           // (terminated)
		.almost_full_data  (),                                                                               // (terminated)
		.almost_empty_data (),                                                                               // (terminated)
		.in_empty          (1'b0),                                                                           // (terminated)
		.out_empty         (),                                                                               // (terminated)
		.in_error          (1'b0),                                                                           // (terminated)
		.out_error         (),                                                                               // (terminated)
		.in_channel        (1'b0),                                                                           // (terminated)
		.out_channel       ()                                                                                // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (101),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_SRC_ID_H              (104),
		.PKT_SRC_ID_L              (103),
		.PKT_DEST_ID_H             (106),
		.PKT_DEST_ID_L             (105),
		.PKT_BURSTWRAP_H           (93),
		.PKT_BURSTWRAP_L           (84),
		.PKT_BYTE_CNT_H            (83),
		.PKT_BYTE_CNT_L            (74),
		.PKT_PROTECTION_H          (110),
		.PKT_PROTECTION_L          (108),
		.PKT_RESPONSE_STATUS_H     (116),
		.PKT_RESPONSE_STATUS_L     (115),
		.PKT_BURST_SIZE_H          (96),
		.PKT_BURST_SIZE_L          (94),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (117),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1)
	) hexport_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pcie_hard_ip_0_pcie_core_clk_clk),                                                //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (hexport_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (hexport_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (hexport_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (hexport_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (hexport_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (hexport_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (hexport_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (hexport_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (hexport_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (hexport_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (hexport_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (hexport_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (hexport_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (hexport_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (hexport_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (hexport_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                 //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                 //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                  //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                         //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                           //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                               //                .channel
		.rf_sink_ready           (hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (hexport_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (hexport_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (hexport_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (hexport_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (hexport_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (hexport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (hexport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (hexport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (hexport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (hexport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (hexport_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (118),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pcie_hard_ip_0_pcie_core_clk_clk),                                                //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (hexport_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (hexport_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (hexport_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (hexport_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (hexport_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (hexport_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (63),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (137),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64),
		.PKT_ADDR_H                (103),
		.PKT_ADDR_L                (72),
		.PKT_TRANS_COMPRESSED_READ (104),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.PKT_TRANS_READ            (107),
		.PKT_TRANS_LOCK            (108),
		.PKT_SRC_ID_H              (140),
		.PKT_SRC_ID_L              (139),
		.PKT_DEST_ID_H             (142),
		.PKT_DEST_ID_L             (141),
		.PKT_BURSTWRAP_H           (129),
		.PKT_BURSTWRAP_L           (120),
		.PKT_BYTE_CNT_H            (119),
		.PKT_BYTE_CNT_L            (110),
		.PKT_PROTECTION_H          (146),
		.PKT_PROTECTION_L          (144),
		.PKT_RESPONSE_STATUS_H     (152),
		.PKT_RESPONSE_STATUS_L     (151),
		.PKT_BURST_SIZE_H          (132),
		.PKT_BURST_SIZE_L          (130),
		.ST_CHANNEL_W              (4),
		.ST_DATA_W                 (153),
		.AVS_BURSTCOUNT_W          (10),
		.SUPPRESS_0_BYTEEN_CMD     (0),
		.PREVENT_FIFO_OVERFLOW     (1)
	) pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent (
		.clk                     (pcie_hard_ip_0_pcie_core_clk_clk),                                                        //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                          //       clk_reset.reset
		.m0_address              (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (cmd_xbar_demux_src3_ready),                                                               //              cp.ready
		.cp_valid                (cmd_xbar_demux_src3_valid),                                                               //                .valid
		.cp_data                 (cmd_xbar_demux_src3_data),                                                                //                .data
		.cp_startofpacket        (cmd_xbar_demux_src3_startofpacket),                                                       //                .startofpacket
		.cp_endofpacket          (cmd_xbar_demux_src3_endofpacket),                                                         //                .endofpacket
		.cp_channel              (cmd_xbar_demux_src3_channel),                                                             //                .channel
		.rf_sink_ready           (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_sink_data    (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.rdata_fifo_src_ready    (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data)         //                .data
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (154),
		.FIFO_DEPTH          (9),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pcie_hard_ip_0_pcie_core_clk_clk),                                                        //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                          // clk_reset.reset
		.in_data           (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                   // (terminated)
		.csr_read          (1'b0),                                                                                    // (terminated)
		.csr_write         (1'b0),                                                                                    // (terminated)
		.csr_readdata      (),                                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                    // (terminated)
		.almost_full_data  (),                                                                                        // (terminated)
		.almost_empty_data (),                                                                                        // (terminated)
		.in_empty          (1'b0),                                                                                    // (terminated)
		.out_empty         (),                                                                                        // (terminated)
		.in_error          (1'b0),                                                                                    // (terminated)
		.out_error         (),                                                                                        // (terminated)
		.in_channel        (1'b0),                                                                                    // (terminated)
		.out_channel       ()                                                                                         // (terminated)
	);

	pcihellocore_addr_router addr_router (
		.sink_ready         (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pcie_hard_ip_0_bar0_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pcie_hard_ip_0_pcie_core_clk_clk),                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                           //       src.ready
		.src_valid          (addr_router_src_valid),                                                           //          .valid
		.src_data           (addr_router_src_data),                                                            //          .data
		.src_channel        (addr_router_src_channel),                                                         //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                      //          .endofpacket
	);

	pcihellocore_id_router id_router (
		.sink_ready         (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pcie_hard_ip_0_cra_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pcie_hard_ip_0_pcie_core_clk_clk),                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_src_ready),                                                           //       src.ready
		.src_valid          (id_router_src_valid),                                                           //          .valid
		.src_data           (id_router_src_data),                                                            //          .data
		.src_channel        (id_router_src_channel),                                                         //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                                                   //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                                                      //          .endofpacket
	);

	pcihellocore_id_router id_router_001 (
		.sink_ready         (inport_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (inport_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (inport_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (inport_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (inport_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pcie_hard_ip_0_pcie_core_clk_clk),                                     //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                       // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                                              //       src.ready
		.src_valid          (id_router_001_src_valid),                                              //          .valid
		.src_data           (id_router_001_src_data),                                               //          .data
		.src_channel        (id_router_001_src_channel),                                            //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                                      //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                                         //          .endofpacket
	);

	pcihellocore_id_router id_router_002 (
		.sink_ready         (hexport_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (hexport_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (hexport_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (hexport_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hexport_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pcie_hard_ip_0_pcie_core_clk_clk),                                      //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                               //       src.ready
		.src_valid          (id_router_002_src_valid),                                               //          .valid
		.src_data           (id_router_002_src_data),                                                //          .data
		.src_channel        (id_router_002_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                          //          .endofpacket
	);

	pcihellocore_id_router_003 id_router_003 (
		.sink_ready         (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (pcie_hard_ip_0_txs_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pcie_hard_ip_0_pcie_core_clk_clk),                                              //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                       //       src.ready
		.src_valid          (id_router_003_src_valid),                                                       //          .valid
		.src_data           (id_router_003_src_data),                                                        //          .data
		.src_channel        (id_router_003_src_channel),                                                     //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                               //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                                  //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (142),
		.PKT_DEST_ID_L             (141),
		.PKT_TRANS_POSTED          (105),
		.PKT_TRANS_WRITE           (106),
		.MAX_OUTSTANDING_RESPONSES (8),
		.PIPELINED                 (0),
		.ST_DATA_W                 (153),
		.ST_CHANNEL_W              (4),
		.VALID_WIDTH               (4),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (119),
		.PKT_BYTE_CNT_L            (110),
		.PKT_BYTEEN_H              (71),
		.PKT_BYTEEN_L              (64)
	) limiter (
		.clk                    (pcie_hard_ip_0_pcie_core_clk_clk), //       clk.clk
		.reset                  (rst_controller_reset_out_reset),   // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),            //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),            //          .valid
		.cmd_sink_data          (addr_router_src_data),             //          .data
		.cmd_sink_channel       (addr_router_src_channel),          //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),    //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),      //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),            //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),             //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),          //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),    //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),      //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),           //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),           //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),         //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),            //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket),   //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),     //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),            //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),            //          .valid
		.rsp_src_data           (limiter_rsp_src_data),             //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),          //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),    //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),      //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)            // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (101),
		.PKT_BYTE_CNT_H            (83),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (96),
		.PKT_BURST_SIZE_L          (94),
		.PKT_BURST_TYPE_H          (98),
		.PKT_BURST_TYPE_L          (97),
		.PKT_BURSTWRAP_H           (93),
		.PKT_BURSTWRAP_L           (84),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (117),
		.ST_CHANNEL_W              (4),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (93),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (1023),
		.BURSTWRAP_CONST_VALUE     (1023)
	) burst_adapter (
		.clk                   (pcie_hard_ip_0_pcie_core_clk_clk),    //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (width_adapter_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_src_data),              //          .data
		.sink0_channel         (width_adapter_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_src_ready),             //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (101),
		.PKT_BYTE_CNT_H            (83),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (96),
		.PKT_BURST_SIZE_L          (94),
		.PKT_BURST_TYPE_H          (98),
		.PKT_BURST_TYPE_L          (97),
		.PKT_BURSTWRAP_H           (93),
		.PKT_BURSTWRAP_L           (84),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (117),
		.ST_CHANNEL_W              (4),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (93),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (1023),
		.BURSTWRAP_CONST_VALUE     (1023)
	) burst_adapter_001 (
		.clk                   (pcie_hard_ip_0_pcie_core_clk_clk),        //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_002_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_002_src_data),              //          .data
		.sink0_channel         (width_adapter_002_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_002_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_002_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_002_src_ready),             //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (101),
		.PKT_BYTE_CNT_H            (83),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (96),
		.PKT_BURST_SIZE_L          (94),
		.PKT_BURST_TYPE_H          (98),
		.PKT_BURST_TYPE_L          (97),
		.PKT_BURSTWRAP_H           (93),
		.PKT_BURSTWRAP_L           (84),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (0),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (117),
		.ST_CHANNEL_W              (4),
		.OUT_BYTE_CNT_H            (76),
		.OUT_BURSTWRAP_H           (93),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (0),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (1023),
		.BURSTWRAP_CONST_VALUE     (1023)
	) burst_adapter_002 (
		.clk                   (pcie_hard_ip_0_pcie_core_clk_clk),        //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (width_adapter_004_src_valid),             //     sink0.valid
		.sink0_data            (width_adapter_004_src_data),              //          .data
		.sink0_channel         (width_adapter_004_src_channel),           //          .channel
		.sink0_startofpacket   (width_adapter_004_src_startofpacket),     //          .startofpacket
		.sink0_endofpacket     (width_adapter_004_src_endofpacket),       //          .endofpacket
		.sink0_ready           (width_adapter_004_src_ready),             //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2)
	) rst_controller (
		.reset_in0  (~pcie_hard_ip_0_pcie_core_reset_reset), // reset_in0.reset
		.clk        (pcie_hard_ip_0_pcie_core_clk_clk),      //       clk.clk
		.reset_out  (rst_controller_reset_out_reset),        // reset_out.reset
		.reset_in1  (1'b0),                                  // (terminated)
		.reset_in2  (1'b0),                                  // (terminated)
		.reset_in3  (1'b0),                                  // (terminated)
		.reset_in4  (1'b0),                                  // (terminated)
		.reset_in5  (1'b0),                                  // (terminated)
		.reset_in6  (1'b0),                                  // (terminated)
		.reset_in7  (1'b0),                                  // (terminated)
		.reset_in8  (1'b0),                                  // (terminated)
		.reset_in9  (1'b0),                                  // (terminated)
		.reset_in10 (1'b0),                                  // (terminated)
		.reset_in11 (1'b0),                                  // (terminated)
		.reset_in12 (1'b0),                                  // (terminated)
		.reset_in13 (1'b0),                                  // (terminated)
		.reset_in14 (1'b0),                                  // (terminated)
		.reset_in15 (1'b0)                                   // (terminated)
	);

	pcihellocore_cmd_xbar_demux cmd_xbar_demux (
		.clk                (pcie_hard_ip_0_pcie_core_clk_clk),  //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_src3_endofpacket)    //           .endofpacket
	);

	pcihellocore_rsp_xbar_demux rsp_xbar_demux (
		.clk                (pcie_hard_ip_0_pcie_core_clk_clk),    //       clk.clk
		.reset              (rst_controller_reset_out_reset),      // clk_reset.reset
		.sink_ready         (width_adapter_001_src_ready),         //      sink.ready
		.sink_channel       (width_adapter_001_src_channel),       //          .channel
		.sink_data          (width_adapter_001_src_data),          //          .data
		.sink_startofpacket (width_adapter_001_src_startofpacket), //          .startofpacket
		.sink_endofpacket   (width_adapter_001_src_endofpacket),   //          .endofpacket
		.sink_valid         (width_adapter_001_src_valid),         //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),           //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),           //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),            //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),         //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),   //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)      //          .endofpacket
	);

	pcihellocore_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (pcie_hard_ip_0_pcie_core_clk_clk),      //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_003_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_003_src_channel),         //          .channel
		.sink_data          (width_adapter_003_src_data),            //          .data
		.sink_startofpacket (width_adapter_003_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_003_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_003_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	pcihellocore_rsp_xbar_demux rsp_xbar_demux_002 (
		.clk                (pcie_hard_ip_0_pcie_core_clk_clk),      //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (width_adapter_005_src_ready),           //      sink.ready
		.sink_channel       (width_adapter_005_src_channel),         //          .channel
		.sink_data          (width_adapter_005_src_data),            //          .data
		.sink_startofpacket (width_adapter_005_src_startofpacket),   //          .startofpacket
		.sink_endofpacket   (width_adapter_005_src_endofpacket),     //          .endofpacket
		.sink_valid         (width_adapter_005_src_valid),           //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	pcihellocore_rsp_xbar_demux rsp_xbar_demux_003 (
		.clk                (pcie_hard_ip_0_pcie_core_clk_clk),      //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	pcihellocore_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (pcie_hard_ip_0_pcie_core_clk_clk),      //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_002_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_003_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (119),
		.IN_PKT_BYTE_CNT_L             (110),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (129),
		.IN_PKT_BURSTWRAP_L            (120),
		.IN_PKT_BURST_SIZE_H           (132),
		.IN_PKT_BURST_SIZE_L           (130),
		.IN_PKT_RESPONSE_STATUS_H      (152),
		.IN_PKT_RESPONSE_STATUS_L      (151),
		.IN_PKT_TRANS_EXCLUSIVE        (109),
		.IN_PKT_BURST_TYPE_H           (134),
		.IN_PKT_BURST_TYPE_L           (133),
		.IN_ST_DATA_W                  (153),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (83),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (96),
		.OUT_PKT_BURST_SIZE_L          (94),
		.OUT_PKT_RESPONSE_STATUS_H     (116),
		.OUT_PKT_RESPONSE_STATUS_L     (115),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (98),
		.OUT_PKT_BURST_TYPE_L          (97),
		.OUT_ST_DATA_W                 (117),
		.ST_CHANNEL_W                  (4),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter (
		.clk                  (pcie_hard_ip_0_pcie_core_clk_clk),  //       clk.clk
		.reset                (rst_controller_reset_out_reset),    // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src0_valid),         //      sink.valid
		.in_channel           (cmd_xbar_demux_src0_channel),       //          .channel
		.in_startofpacket     (cmd_xbar_demux_src0_startofpacket), //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src0_endofpacket),   //          .endofpacket
		.in_ready             (cmd_xbar_demux_src0_ready),         //          .ready
		.in_data              (cmd_xbar_demux_src0_data),          //          .data
		.out_endofpacket      (width_adapter_src_endofpacket),     //       src.endofpacket
		.out_data             (width_adapter_src_data),            //          .data
		.out_channel          (width_adapter_src_channel),         //          .channel
		.out_valid            (width_adapter_src_valid),           //          .valid
		.out_ready            (width_adapter_src_ready),           //          .ready
		.out_startofpacket    (width_adapter_src_startofpacket),   //          .startofpacket
		.in_command_size_data (3'b000)                             // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (83),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (93),
		.IN_PKT_BURSTWRAP_L            (84),
		.IN_PKT_BURST_SIZE_H           (96),
		.IN_PKT_BURST_SIZE_L           (94),
		.IN_PKT_RESPONSE_STATUS_H      (116),
		.IN_PKT_RESPONSE_STATUS_L      (115),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (98),
		.IN_PKT_BURST_TYPE_L           (97),
		.IN_ST_DATA_W                  (117),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (119),
		.OUT_PKT_BYTE_CNT_L            (110),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_PKT_BURST_SIZE_H          (132),
		.OUT_PKT_BURST_SIZE_L          (130),
		.OUT_PKT_RESPONSE_STATUS_H     (152),
		.OUT_PKT_RESPONSE_STATUS_L     (151),
		.OUT_PKT_TRANS_EXCLUSIVE       (109),
		.OUT_PKT_BURST_TYPE_H          (134),
		.OUT_PKT_BURST_TYPE_L          (133),
		.OUT_ST_DATA_W                 (153),
		.ST_CHANNEL_W                  (4),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_001 (
		.clk                  (pcie_hard_ip_0_pcie_core_clk_clk),    //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_src_valid),                 //      sink.valid
		.in_channel           (id_router_src_channel),               //          .channel
		.in_startofpacket     (id_router_src_startofpacket),         //          .startofpacket
		.in_endofpacket       (id_router_src_endofpacket),           //          .endofpacket
		.in_ready             (id_router_src_ready),                 //          .ready
		.in_data              (id_router_src_data),                  //          .data
		.out_endofpacket      (width_adapter_001_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_001_src_data),          //          .data
		.out_channel          (width_adapter_001_src_channel),       //          .channel
		.out_valid            (width_adapter_001_src_valid),         //          .valid
		.out_ready            (width_adapter_001_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_001_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (119),
		.IN_PKT_BYTE_CNT_L             (110),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (129),
		.IN_PKT_BURSTWRAP_L            (120),
		.IN_PKT_BURST_SIZE_H           (132),
		.IN_PKT_BURST_SIZE_L           (130),
		.IN_PKT_RESPONSE_STATUS_H      (152),
		.IN_PKT_RESPONSE_STATUS_L      (151),
		.IN_PKT_TRANS_EXCLUSIVE        (109),
		.IN_PKT_BURST_TYPE_H           (134),
		.IN_PKT_BURST_TYPE_L           (133),
		.IN_ST_DATA_W                  (153),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (83),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (96),
		.OUT_PKT_BURST_SIZE_L          (94),
		.OUT_PKT_RESPONSE_STATUS_H     (116),
		.OUT_PKT_RESPONSE_STATUS_L     (115),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (98),
		.OUT_PKT_BURST_TYPE_L          (97),
		.OUT_ST_DATA_W                 (117),
		.ST_CHANNEL_W                  (4),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_002 (
		.clk                  (pcie_hard_ip_0_pcie_core_clk_clk),    //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src1_valid),           //      sink.valid
		.in_channel           (cmd_xbar_demux_src1_channel),         //          .channel
		.in_startofpacket     (cmd_xbar_demux_src1_startofpacket),   //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src1_endofpacket),     //          .endofpacket
		.in_ready             (cmd_xbar_demux_src1_ready),           //          .ready
		.in_data              (cmd_xbar_demux_src1_data),            //          .data
		.out_endofpacket      (width_adapter_002_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_002_src_data),          //          .data
		.out_channel          (width_adapter_002_src_channel),       //          .channel
		.out_valid            (width_adapter_002_src_valid),         //          .valid
		.out_ready            (width_adapter_002_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_002_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (83),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (93),
		.IN_PKT_BURSTWRAP_L            (84),
		.IN_PKT_BURST_SIZE_H           (96),
		.IN_PKT_BURST_SIZE_L           (94),
		.IN_PKT_RESPONSE_STATUS_H      (116),
		.IN_PKT_RESPONSE_STATUS_L      (115),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (98),
		.IN_PKT_BURST_TYPE_L           (97),
		.IN_ST_DATA_W                  (117),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (119),
		.OUT_PKT_BYTE_CNT_L            (110),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_PKT_BURST_SIZE_H          (132),
		.OUT_PKT_BURST_SIZE_L          (130),
		.OUT_PKT_RESPONSE_STATUS_H     (152),
		.OUT_PKT_RESPONSE_STATUS_L     (151),
		.OUT_PKT_TRANS_EXCLUSIVE       (109),
		.OUT_PKT_BURST_TYPE_H          (134),
		.OUT_PKT_BURST_TYPE_L          (133),
		.OUT_ST_DATA_W                 (153),
		.ST_CHANNEL_W                  (4),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_003 (
		.clk                  (pcie_hard_ip_0_pcie_core_clk_clk),    //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_001_src_valid),             //      sink.valid
		.in_channel           (id_router_001_src_channel),           //          .channel
		.in_startofpacket     (id_router_001_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_001_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_001_src_ready),             //          .ready
		.in_data              (id_router_001_src_data),              //          .data
		.out_endofpacket      (width_adapter_003_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_003_src_data),          //          .data
		.out_channel          (width_adapter_003_src_channel),       //          .channel
		.out_valid            (width_adapter_003_src_valid),         //          .valid
		.out_ready            (width_adapter_003_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_003_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (103),
		.IN_PKT_ADDR_L                 (72),
		.IN_PKT_DATA_H                 (63),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (71),
		.IN_PKT_BYTEEN_L               (64),
		.IN_PKT_BYTE_CNT_H             (119),
		.IN_PKT_BYTE_CNT_L             (110),
		.IN_PKT_TRANS_COMPRESSED_READ  (104),
		.IN_PKT_BURSTWRAP_H            (129),
		.IN_PKT_BURSTWRAP_L            (120),
		.IN_PKT_BURST_SIZE_H           (132),
		.IN_PKT_BURST_SIZE_L           (130),
		.IN_PKT_RESPONSE_STATUS_H      (152),
		.IN_PKT_RESPONSE_STATUS_L      (151),
		.IN_PKT_TRANS_EXCLUSIVE        (109),
		.IN_PKT_BURST_TYPE_H           (134),
		.IN_PKT_BURST_TYPE_L           (133),
		.IN_ST_DATA_W                  (153),
		.OUT_PKT_ADDR_H                (67),
		.OUT_PKT_ADDR_L                (36),
		.OUT_PKT_DATA_H                (31),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (35),
		.OUT_PKT_BYTEEN_L              (32),
		.OUT_PKT_BYTE_CNT_H            (83),
		.OUT_PKT_BYTE_CNT_L            (74),
		.OUT_PKT_TRANS_COMPRESSED_READ (68),
		.OUT_PKT_BURST_SIZE_H          (96),
		.OUT_PKT_BURST_SIZE_L          (94),
		.OUT_PKT_RESPONSE_STATUS_H     (116),
		.OUT_PKT_RESPONSE_STATUS_L     (115),
		.OUT_PKT_TRANS_EXCLUSIVE       (73),
		.OUT_PKT_BURST_TYPE_H          (98),
		.OUT_PKT_BURST_TYPE_L          (97),
		.OUT_ST_DATA_W                 (117),
		.ST_CHANNEL_W                  (4),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_004 (
		.clk                  (pcie_hard_ip_0_pcie_core_clk_clk),    //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (cmd_xbar_demux_src2_valid),           //      sink.valid
		.in_channel           (cmd_xbar_demux_src2_channel),         //          .channel
		.in_startofpacket     (cmd_xbar_demux_src2_startofpacket),   //          .startofpacket
		.in_endofpacket       (cmd_xbar_demux_src2_endofpacket),     //          .endofpacket
		.in_ready             (cmd_xbar_demux_src2_ready),           //          .ready
		.in_data              (cmd_xbar_demux_src2_data),            //          .data
		.out_endofpacket      (width_adapter_004_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_004_src_data),          //          .data
		.out_channel          (width_adapter_004_src_channel),       //          .channel
		.out_valid            (width_adapter_004_src_valid),         //          .valid
		.out_ready            (width_adapter_004_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_004_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	altera_merlin_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (83),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (93),
		.IN_PKT_BURSTWRAP_L            (84),
		.IN_PKT_BURST_SIZE_H           (96),
		.IN_PKT_BURST_SIZE_L           (94),
		.IN_PKT_RESPONSE_STATUS_H      (116),
		.IN_PKT_RESPONSE_STATUS_L      (115),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (98),
		.IN_PKT_BURST_TYPE_L           (97),
		.IN_ST_DATA_W                  (117),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (119),
		.OUT_PKT_BYTE_CNT_L            (110),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_PKT_BURST_SIZE_H          (132),
		.OUT_PKT_BURST_SIZE_L          (130),
		.OUT_PKT_RESPONSE_STATUS_H     (152),
		.OUT_PKT_RESPONSE_STATUS_L     (151),
		.OUT_PKT_TRANS_EXCLUSIVE       (109),
		.OUT_PKT_BURST_TYPE_H          (134),
		.OUT_PKT_BURST_TYPE_L          (133),
		.OUT_ST_DATA_W                 (153),
		.ST_CHANNEL_W                  (4),
		.OPTIMIZE_FOR_RSP              (0)
	) width_adapter_005 (
		.clk                  (pcie_hard_ip_0_pcie_core_clk_clk),    //       clk.clk
		.reset                (rst_controller_reset_out_reset),      // clk_reset.reset
		.in_valid             (id_router_002_src_valid),             //      sink.valid
		.in_channel           (id_router_002_src_channel),           //          .channel
		.in_startofpacket     (id_router_002_src_startofpacket),     //          .startofpacket
		.in_endofpacket       (id_router_002_src_endofpacket),       //          .endofpacket
		.in_ready             (id_router_002_src_ready),             //          .ready
		.in_data              (id_router_002_src_data),              //          .data
		.out_endofpacket      (width_adapter_005_src_endofpacket),   //       src.endofpacket
		.out_data             (width_adapter_005_src_data),          //          .data
		.out_channel          (width_adapter_005_src_channel),       //          .channel
		.out_valid            (width_adapter_005_src_valid),         //          .valid
		.out_ready            (width_adapter_005_src_ready),         //          .ready
		.out_startofpacket    (width_adapter_005_src_startofpacket), //          .startofpacket
		.in_command_size_data (3'b000)                               // (terminated)
	);

	pcihellocore_irq_mapper irq_mapper (
		.clk        (pcie_hard_ip_0_pcie_core_clk_clk),      //       clk.clk
		.reset      (~pcie_hard_ip_0_pcie_core_reset_reset), // clk_reset.reset
		.sender_irq (irq_synchronizer_receiver_irq)          //    sender.irq
	);

	altera_irq_clock_crosser #(
		.IRQ_WIDTH (16)
	) irq_synchronizer (
		.receiver_clk   (pcie_hard_ip_0_pcie_core_clk_clk),      //       receiver_clk.clk
		.sender_clk     (pcie_hard_ip_0_pcie_core_clk_clk),      //         sender_clk.clk
		.receiver_reset (~pcie_hard_ip_0_pcie_core_reset_reset), // receiver_clk_reset.reset
		.sender_reset   (~pcie_hard_ip_0_pcie_core_reset_reset), //   sender_clk_reset.reset
		.receiver_irq   (irq_synchronizer_receiver_irq),         //           receiver.irq
		.sender_irq     (pcie_hard_ip_0_rxm_irq_irq)             //             sender.irq
	);

endmodule
